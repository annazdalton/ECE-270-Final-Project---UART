//will add parity check logic
module parityChecker(
    input logic [7:0] sipo_i,
    input logic parity_en, parity_bit, //parity_bit is data_i from transmitter
    output logic parity_error
);

endmodule
