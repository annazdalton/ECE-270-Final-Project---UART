module transmitter_parityGen();

endmodule