module transmitterMux(
    input logic [7:0] data_i,
    input logic shift_en,
    output logic piso_o
);


endmodule 